module pop_count(g, c, a)
input a, c, g
