module pop_count()
